05 06 2018
12 00 00
350
Place
Description
4
DDDD
DDD
DD
D
06 04 2018
10 00 00
350
Ivano-Frankivsk
Sightseeing
2
Bodia
Dima
12 05 2019
23 00 00
120
Lviv
Night walk
4
Lisa
Nastia
Bodia
Nazar
12 00 00
12 00 00
32
Place
DDDDDDD
3
One
Two
Three
12 02 2019
12:00:00
120

Des
2
Dime
Nino
